`timescale 1 ns / 1 ps

/*

MPS AXI4_Lite_S01 Module
개발 4팀 전경원 차장

24.06.10 :	최초 생성
24.07.08 :	DPBRAM Test용 AXI 추가
			직병렬 기능 추가 및 업데이트에 따라서 slv_reg 주소 변경할 수도 있음

			Name					slv_reg
			o_test_dpbram_addr : 	62
			o_test_dpbram_en : 		63[0]
			o_test_dpbram_w_en : 	63[1]
			o_test_dpbram_wdata : 	50
			i_test_dpbram_rdata : 	7

이성진 차장의 퇴사로 인하여 MPS PL 프로그래밍

- 안쓰는 Reg 정리 필요

REG에 쓰는게 input (PL -> PS)
REG를 읽는게 output (PS -> PL)
input 주석처리

*/

module AXI4_Lite_S01 #
(
	parameter integer C_S_AXI_DATA_WIDTH	= 0,
	parameter integer C_S_AXI_ADDR_WIDTH	= 0
)
(
	//Write
	output reg [31:0] 		o_c_factor,
	output reg [31:0] 		o_v_factor,
	output reg 	[31:0]		o_WF_total_count,
	output reg 				o_WF_BRAM_WE,
	output reg 				o_WF_start_count,
	output reg 				o_WF_reset_count,
	output reg 				o_WF_mode_sel,
	output reg 	[9:0]		o_WF_addr,
	output reg 	[31:0]		o_WF_data,
	output reg 	[15:0]		o_WF_dsp,
	output reg 				o_Ready,
	output reg 				o_Hart_beat,
	output reg 	[15:0]		o_Write_Index,
	output reg 	[31:0]		o_Write_DATA,

	output reg [9:0]		o_test_dpbram_addr,		// Test용 DPBRAM ADDR
	output reg 				o_test_dpbram_en,		// Test용 DPBRAM Enable
	output reg 				o_test_dpbram_w_en,		// Test용 DPBRAM Wirte Flag
	output reg 				o_test_dpbram_DSP_intr,	// Test용 DPBRAM DSP Interrupt
	output reg [15:0]		o_test_dpbram_wdata,	// Test용 DPBRAM Write Data

	//Read
	input 					i_WF_INT_0,
	input 					i_WF_INT_500,
	input [31:0]			i_WF_current_count,
	input 					i_valid,
	input 					i_DSP_fail,
	input 					i_DSP_nENPWM,
	input [31:0]			i_Float_ADC_C,
	input [31:0]			i_Float_ADC_V,
	input [31:0]			i_DSP_Duty,
	input [15:0]			i_DSP_FaultNum,
	input [31:0]			i_DSP_System_Status,
	input [15:0]			i_DSP_EIS,
	input [31:0]			i_DSP_RLoad,
	input [15:0]			i_DSP_MPS_TYPE,
	input [31:0]			i_DSP_SetCurrRD,
	input [31:0]			i_DSP_DEGCurrentRD,
	input [31:0]			i_DSP_DEGPeriod,
	input [31:0]			i_DSP_OverCurrent,
	input [31:0]			i_DSP_LowVoltage,
	input [31:0]			i_DSP_OverVoltage,
	input [31:0]			i_DSP_OverTemp,
	input [31:0]			i_DSP_CurrentHighLimit,
	input [31:0]			i_DSP_Vpgain,
	input [31:0]			i_DSP_ViGain,
	input [31:0]			i_DSP_CurrentPgain,
	input [31:0]			i_DSP_CurrentIgain,
	input [31:0]			i_DSP_Max_Duty,
	input [15:0]			i_DSP_DSP_Code,
	input [15:0]			i_DSP_SlewRate,
	input [15:0]			i_DSP_osc_state,
	input [15:0]			i_DSP_remote_state,
	input [31:0]			i_DSP_regulation_time,
	input [31:0]			i_DSP_Current_Factor,
	input [31:0]			i_DSP_Voltage_Factor,
	input [31:0]			i_DSP_Input_Voltage_Factor,
	input [31:0]			i_DSP_Current_Offset_Set,
	input [15:0]			i_DSP_Deadband_Set,
	input [15:0]			i_DSP_Dual_Offset_Deadband_Set,
	input [31:0]			i_DSP_PI_Max_V,
	input [31:0]			i_DSP_PI_Min_V,
	input [31:0]			i_DSP_Eruption_V,
	input [31:0]			i_DSP_Eruption_C,
	input [31:0]			i_F_DSP_ADC_C,
	input [31:0]			i_F_DSP_ADC_V,

	input [15:0]			i_test_dpbram_rdata,		// Test용 DPBRAM Read Data


	// User ports ends
	// Do not modify the ports beyond this line
	// Global Clock Signal
	input wire  S_AXI_ACLK,
	// Global Reset Signal. This Signal is Active LOW
	input wire  S_AXI_ARESETN,
	// Write address (issued by master, acceped by Slave)
	input wire [C_S_AXI_ADDR_WIDTH-1 : 0] S_AXI_AWADDR,
	// Write channel Protection type. This signal indicates the
		// privilege and security level of the transaction, and whether
		// the transaction is a data access or an instruction access.
	input wire [2 : 0] S_AXI_AWPROT,
	// Write address valid. This signal indicates that the master signaling
		// valid write address and control information.
	input wire  S_AXI_AWVALID,
	// Write address ready. This signal indicates that the slave is ready
		// to accept an address and associated control signals.
	output wire  S_AXI_AWREADY,
	// Write data (issued by master, acceped by Slave) 
	input wire [C_S_AXI_DATA_WIDTH-1 : 0] S_AXI_WDATA,
	// Write strobes. This signal indicates which byte lanes hold
		// valid data. There is one write strobe bit for each eight
		// bits of the write data bus.    
	input wire [(C_S_AXI_DATA_WIDTH/8)-1 : 0] S_AXI_WSTRB,
	// Write valid. This signal indicates that valid write
		// data and strobes are available.
	input wire  S_AXI_WVALID,
	// Write ready. This signal indicates that the slave
		// can accept the write data.
	output wire  S_AXI_WREADY,
	// Write response. This signal indicates the status
		// of the write transaction.
	output wire [1 : 0] S_AXI_BRESP,
	// Write response valid. This signal indicates that the channel
		// is signaling a valid write response.
	output wire  S_AXI_BVALID,
	// Response ready. This signal indicates that the master
		// can accept a write response.
	input wire  S_AXI_BREADY,
	// Read address (issued by master, acceped by Slave)
	input wire [C_S_AXI_ADDR_WIDTH-1 : 0] S_AXI_ARADDR,
	// Protection type. This signal indicates the privilege
		// and security level of the transaction, and whether the
		// transaction is a data access or an instruction access.
	input wire [2 : 0] S_AXI_ARPROT,
	// Read address valid. This signal indicates that the channel
		// is signaling valid read address and control information.
	input wire  S_AXI_ARVALID,
	// Read address ready. This signal indicates that the slave is
		// ready to accept an address and associated control signals.
	output wire  S_AXI_ARREADY,
	// Read data (issued by slave)
	output wire [C_S_AXI_DATA_WIDTH-1 : 0] S_AXI_RDATA,
	// Read response. This signal indicates the status of the
		// read transfer.
	output wire [1 : 0] S_AXI_RRESP,
	// Read valid. This signal indicates that the channel is
		// signaling the required read data.
	output wire  S_AXI_RVALID,
	// Read ready. This signal indicates that the master can
		// accept the read data and response information.
	input wire  S_AXI_RREADY
);

	// AXI4LITE signals
	reg [C_S_AXI_ADDR_WIDTH-1 : 0] 	axi_awaddr;
	reg  	axi_awready;
	reg  	axi_wready;
	reg [1 : 0] 	axi_bresp;
	reg  	axi_bvalid;
	reg [C_S_AXI_ADDR_WIDTH-1 : 0] 	axi_araddr;
	reg  	axi_arready;
	reg [C_S_AXI_DATA_WIDTH-1 : 0] 	axi_rdata;
	reg [1 : 0] 	axi_rresp;
	reg  	axi_rvalid;

	// Example-specific design signals
	// local parameter for addressing 32 bit / 64 bit C_S_AXI_DATA_WIDTH
	// ADDR_LSB is used for addressing 32/64 bit registers/memories
	// ADDR_LSB = 2 for 32 bits (n downto 2)
	// ADDR_LSB = 3 for 64 bits (n downto 3)
	localparam integer ADDR_LSB = (C_S_AXI_DATA_WIDTH/32) + 1;
	localparam integer OPT_MEM_ADDR_BITS = 5;
	//----------------------------------------------
	//-- Signals for user logic register space example
	//------------------------------------------------
	//-- Number of Slave Registers 64
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg0;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg1;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg2;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg3;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg4;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg5;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg6;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg7;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg8;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg9;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg10;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg11;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg12;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg13;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg14;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg15;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg16;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg17;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg18;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg19;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg20;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg21;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg22;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg23;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg24;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg25;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg26;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg27;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg28;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg29;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg30;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg31;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg32;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg33;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg34;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg35;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg36;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg37;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg38;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg39;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg40;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg41;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg42;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg43;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg44;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg45;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg46;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg47;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg48;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg49;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg50;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg51;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg52;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg53;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg54;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg55;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg56;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg57;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg58;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg59;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg60;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg61;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg62;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg63;

	wire	 slv_reg_rden;
	wire	 slv_reg_wren;
	reg [C_S_AXI_DATA_WIDTH-1:0]	 reg_data_out;
	integer	 byte_index;
	reg	 aw_en;

	// I/O Connections assignments

	assign S_AXI_AWREADY	= axi_awready;
	assign S_AXI_WREADY	= axi_wready;
	assign S_AXI_BRESP	= axi_bresp;
	assign S_AXI_BVALID	= axi_bvalid;
	assign S_AXI_ARREADY	= axi_arready;
	assign S_AXI_RDATA	= axi_rdata;
	assign S_AXI_RRESP	= axi_rresp;
	assign S_AXI_RVALID	= axi_rvalid;
	// Implement axi_awready generation
	// axi_awready is asserted for one S_AXI_ACLK clock cycle when both
	// S_AXI_AWVALID and S_AXI_WVALID are asserted. axi_awready is
	// de-asserted when reset is low.

	always @( posedge S_AXI_ACLK )
	begin
	  if ( S_AXI_ARESETN == 1'b0 )
	    begin
	      axi_awready <= 1'b0;
	      aw_en <= 1'b1;
	    end 
	  else
	    begin    
	      if (~axi_awready && S_AXI_AWVALID && S_AXI_WVALID && aw_en)
	        begin
	          // slave is ready to accept write address when 
	          // there is a valid write address and write data
	          // on the write address and data bus. This design 
	          // expects no outstanding transactions. 
	          axi_awready <= 1'b1;
	          aw_en <= 1'b0;
	        end
	        else if (S_AXI_BREADY && axi_bvalid)
	            begin
	              aw_en <= 1'b1;
	              axi_awready <= 1'b0;
	            end
	      else           
	        begin
	          axi_awready <= 1'b0;
	        end
	    end 
	end       

	// Implement axi_awaddr latching
	// This process is used to latch the address when both 
	// S_AXI_AWVALID and S_AXI_WVALID are valid. 

	always @( posedge S_AXI_ACLK )
	begin
	  if ( S_AXI_ARESETN == 1'b0 )
	    begin
	      axi_awaddr <= 0;
	    end 
	  else
	    begin    
	      if (~axi_awready && S_AXI_AWVALID && S_AXI_WVALID && aw_en)
	        begin
	          // Write Address latching 
	          axi_awaddr <= S_AXI_AWADDR;
	        end
	    end 
	end       

	// Implement axi_wready generation
	// axi_wready is asserted for one S_AXI_ACLK clock cycle when both
	// S_AXI_AWVALID and S_AXI_WVALID are asserted. axi_wready is 
	// de-asserted when reset is low. 

	always @( posedge S_AXI_ACLK )
	begin
	  if ( S_AXI_ARESETN == 1'b0 )
	    begin
	      axi_wready <= 1'b0;
	    end 
	  else
	    begin    
	      if (~axi_wready && S_AXI_WVALID && S_AXI_AWVALID && aw_en )
	        begin
	          // slave is ready to accept write data when 
	          // there is a valid write address and write data
	          // on the write address and data bus. This design 
	          // expects no outstanding transactions. 
	          axi_wready <= 1'b1;
	        end
	      else
	        begin
	          axi_wready <= 1'b0;
	        end
	    end 
	end       

	// Implement memory mapped register select and write logic generation
	// The write data is accepted and written to memory mapped registers when
	// axi_awready, S_AXI_WVALID, axi_wready and S_AXI_WVALID are asserted. Write strobes are used to
	// select byte enables of slave registers while writing.
	// These registers are cleared when reset (active low) is applied.
	// Slave register write enable is asserted when valid address and data are available
	// and the slave is ready to accept the write address and write data.
	assign slv_reg_wren = axi_wready && S_AXI_WVALID && axi_awready && S_AXI_AWVALID;

	always @( posedge S_AXI_ACLK )
	begin
	  if ( S_AXI_ARESETN == 1'b0 )
	    begin
	      slv_reg0 <= 0;
	    //   slv_reg1 <= 0;
	    //   slv_reg2 <= 0;
	      slv_reg3 <= 0;
	      slv_reg4 <= 0;
	      slv_reg5 <= 0;
	      slv_reg6 <= 0;
	    //   slv_reg7 <= 0;
	      slv_reg8 <= 0;
	      slv_reg9 <= 0;
	    //   slv_reg10 <= 0;
	    //   slv_reg11 <= 0;
	      slv_reg12 <= 0;
	    //   slv_reg13 <= 0;
	      slv_reg14 <= 0;
	      slv_reg15 <= 0;
	    //   slv_reg16 <= 0;
	    //   slv_reg17 <= 0;
	    //   slv_reg18 <= 0;
	    //   slv_reg19 <= 0;
	    //   slv_reg20 <= 0;
	    //   slv_reg21 <= 0;
	    //   slv_reg22 <= 0;
	    //   slv_reg23 <= 0;
	    //   slv_reg24 <= 0;
	    //   slv_reg25 <= 0;
	    //   slv_reg26 <= 0;
	    //   slv_reg27 <= 0;
	    //   slv_reg28 <= 0;
	    //   slv_reg29 <= 0;
	    //   slv_reg30 <= 0;
	    //   slv_reg31 <= 0;
	    //   slv_reg32 <= 0;
	    //   slv_reg33 <= 0;
	    //   slv_reg34 <= 0;
	    //   slv_reg35 <= 0;
	    //   slv_reg36 <= 0;
	    //   slv_reg37 <= 0;
	    //   slv_reg38 <= 0;
	    //   slv_reg39 <= 0;
	    //   slv_reg40 <= 0;
	    //   slv_reg41 <= 0;
	    //   slv_reg42 <= 0;
	    //   slv_reg43 <= 0;
	    //   slv_reg44 <= 0;
	    //   slv_reg45 <= 0;
	    //   slv_reg46 <= 0;
	    //   slv_reg47 <= 0;
	    //   slv_reg48 <= 0;
	    //   slv_reg49 <= 0;
	    //   slv_reg50 <= 0;
	    //   slv_reg51 <= 0;
	      slv_reg52 <= 0;
	      slv_reg53 <= 0;
	      slv_reg54 <= 0;
	      slv_reg55 <= 0;
	      slv_reg56 <= 0;
	      slv_reg57 <= 0;
	      slv_reg58 <= 0;
	      slv_reg59 <= 0;
	      slv_reg60 <= 0;
	      slv_reg61 <= 0;
	      slv_reg62 <= 0;
	      slv_reg63 <= 0;
	    end 
	  else begin
	    if (slv_reg_wren)
	      begin
	        case ( axi_awaddr[ADDR_LSB+OPT_MEM_ADDR_BITS:ADDR_LSB] )
	          7'h00:
	            for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	              if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	                // Respective byte enables are asserted as per write strobes 
	                // Slave register 0
	                slv_reg0[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	              end  
	        //   7'h01:
	        //     for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	        //       if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	        //         // Respective byte enables are asserted as per write strobes 
	        //         // Slave register 1
	        //         slv_reg1[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	        //       end  
	        //   7'h02:
	        //     for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	        //       if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	        //         // Respective byte enables are asserted as per write strobes 
	        //         // Slave register 2
	        //         slv_reg2[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	        //       end  
	          7'h03:
	            for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	              if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	                // Respective byte enables are asserted as per write strobes 
	                // Slave register 3
	                slv_reg3[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	              end  
	          7'h04:
	            for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	              if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	                // Respective byte enables are asserted as per write strobes 
	                // Slave register 4
	                slv_reg4[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	              end  
	          7'h05:
	            for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	              if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	                // Respective byte enables are asserted as per write strobes 
	                // Slave register 5
	                slv_reg5[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	              end  
	          7'h06:
	            for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	              if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	                // Respective byte enables are asserted as per write strobes 
	                // Slave register 6
	                slv_reg6[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	              end  
	        //   7'h07:
	        //     for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	        //       if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	        //         // Respective byte enables are asserted as per write strobes 
	        //         // Slave register 7
	        //         slv_reg7[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	        //       end  
	          7'h08:
	            for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	              if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	                // Respective byte enables are asserted as per write strobes 
	                // Slave register 8
	                slv_reg8[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	              end  
	          7'h09:
	            for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	              if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	                // Respective byte enables are asserted as per write strobes 
	                // Slave register 9
	                slv_reg9[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	              end  
	        //   7'h0A:
	        //     for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	        //       if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	        //         // Respective byte enables are asserted as per write strobes 
	        //         // Slave register 10
	        //         slv_reg10[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	        //       end  
	        //   7'h0B:
	        //     for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	        //       if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	        //         // Respective byte enables are asserted as per write strobes 
	        //         // Slave register 11
	        //         slv_reg11[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	        //       end  
	          7'h0C:
	            for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	              if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	                // Respective byte enables are asserted as per write strobes 
	                // Slave register 12
	                slv_reg12[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	              end  
	        //   7'h0D:
	        //     for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	        //       if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	        //         // Respective byte enables are asserted as per write strobes 
	        //         // Slave register 13
	        //         slv_reg13[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	        //       end  
	          7'h0E:
	            for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	              if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	                // Respective byte enables are asserted as per write strobes 
	                // Slave register 14
	                slv_reg14[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	              end  
	          7'h0F:
	            for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	              if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	                // Respective byte enables are asserted as per write strobes 
	                // Slave register 15
	                slv_reg15[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	              end  
	        //   7'h10:
	        //     for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	        //       if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	        //         // Respective byte enables are asserted as per write strobes 
	        //         // Slave register 16
	        //         slv_reg16[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	        //       end  
	        //   7'h11:
	        //     for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	        //       if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	        //         // Respective byte enables are asserted as per write strobes 
	        //         // Slave register 17
	        //         slv_reg17[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	        //       end  
	        //   7'h12:
	        //     for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	        //       if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	        //         // Respective byte enables are asserted as per write strobes 
	        //         // Slave register 18
	        //         slv_reg18[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	        //       end  
	        //   7'h13:
	        //     for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	        //       if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	        //         // Respective byte enables are asserted as per write strobes 
	        //         // Slave register 19
	        //         slv_reg19[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	        //       end  
	        //   7'h14:
	        //     for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	        //       if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	        //         // Respective byte enables are asserted as per write strobes 
	        //         // Slave register 20
	        //         slv_reg20[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	        //       end  
	        //   7'h15:
	        //     for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	        //       if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	        //         // Respective byte enables are asserted as per write strobes 
	        //         // Slave register 21
	        //         slv_reg21[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	        //       end  
	        //   7'h16:
	        //     for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	        //       if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	        //         // Respective byte enables are asserted as per write strobes 
	        //         // Slave register 22
	        //         slv_reg22[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	        //       end  
	        //   7'h17:
	        //     for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	        //       if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	        //         // Respective byte enables are asserted as per write strobes 
	        //         // Slave register 23
	        //         slv_reg23[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	        //       end  
	        //   7'h18:
	        //     for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	        //       if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	        //         // Respective byte enables are asserted as per write strobes 
	        //         // Slave register 24
	        //         slv_reg24[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	        //       end  
	        //   7'h19:
	        //     for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	        //       if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	        //         // Respective byte enables are asserted as per write strobes 
	        //         // Slave register 25
	        //         slv_reg25[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	        //       end  
	        //   7'h1A:
	        //     for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	        //       if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	        //         // Respective byte enables are asserted as per write strobes 
	        //         // Slave register 26
	        //         slv_reg26[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	        //       end  
	        //   7'h1B:
	        //     for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	        //       if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	        //         // Respective byte enables are asserted as per write strobes 
	        //         // Slave register 27
	        //         slv_reg27[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	        //       end  
	        //   7'h1C:
	        //     for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	        //       if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	        //         // Respective byte enables are asserted as per write strobes 
	        //         // Slave register 28
	        //         slv_reg28[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	        //       end  
	        //   7'h1D:
	        //     for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	        //       if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	        //         // Respective byte enables are asserted as per write strobes 
	        //         // Slave register 29
	        //         slv_reg29[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	        //       end  
	        //   7'h1E:
	        //     for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	        //       if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	        //         // Respective byte enables are asserted as per write strobes 
	        //         // Slave register 30
	        //         slv_reg30[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	        //       end  
	        //   7'h1F:
	        //     for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	        //       if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	        //         // Respective byte enables are asserted as per write strobes 
	        //         // Slave register 31
	        //         slv_reg31[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	        //       end  
	        //   7'h20:
	        //     for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	        //       if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	        //         // Respective byte enables are asserted as per write strobes 
	        //         // Slave register 32
	        //         slv_reg32[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	        //       end  
	        //   7'h21:
	        //     for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	        //       if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	        //         // Respective byte enables are asserted as per write strobes 
	        //         // Slave register 33
	        //         slv_reg33[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	        //       end  
	        //   7'h22:
	        //     for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	        //       if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	        //         // Respective byte enables are asserted as per write strobes 
	        //         // Slave register 34
	        //         slv_reg34[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	        //       end  
	        //   7'h23:
	        //     for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	        //       if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	        //         // Respective byte enables are asserted as per write strobes 
	        //         // Slave register 35
	        //         slv_reg35[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	        //       end  
	        //   7'h24:
	        //     for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	        //       if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	        //         // Respective byte enables are asserted as per write strobes 
	        //         // Slave register 36
	        //         slv_reg36[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	        //       end  
	        //   7'h25:
	        //     for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	        //       if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	        //         // Respective byte enables are asserted as per write strobes 
	        //         // Slave register 37
	        //         slv_reg37[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	        //       end  
	        //   7'h26:
	        //     for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	        //       if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	        //         // Respective byte enables are asserted as per write strobes 
	        //         // Slave register 38
	        //         slv_reg38[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	        //       end  
	        //   7'h27:
	        //     for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	        //       if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	        //         // Respective byte enables are asserted as per write strobes 
	        //         // Slave register 39
	        //         slv_reg39[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	        //       end  
	        //   7'h28:
	        //     for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	        //       if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	        //         // Respective byte enables are asserted as per write strobes 
	        //         // Slave register 40
	        //         slv_reg40[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	        //       end  
	        //   7'h29:
	        //     for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	        //       if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	        //         // Respective byte enables are asserted as per write strobes 
	        //         // Slave register 41
	        //         slv_reg41[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	        //       end  
	        //   7'h2A:
	        //     for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	        //       if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	        //         // Respective byte enables are asserted as per write strobes 
	        //         // Slave register 42
	        //         slv_reg42[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	        //       end  
	        //   7'h2B:
	        //     for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	        //       if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	        //         // Respective byte enables are asserted as per write strobes 
	        //         // Slave register 43
	        //         slv_reg43[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	        //       end  
	        //   7'h2C:
	        //     for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	        //       if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	        //         // Respective byte enables are asserted as per write strobes 
	        //         // Slave register 44
	        //         slv_reg44[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	        //       end  
	        //   7'h2D:
	        //     for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	        //       if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	        //         // Respective byte enables are asserted as per write strobes 
	        //         // Slave register 45
	        //         slv_reg45[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	        //       end  
	        //   7'h2E:
	        //     for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	        //       if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	        //         // Respective byte enables are asserted as per write strobes 
	        //         // Slave register 46
	        //         slv_reg46[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	        //       end  
	        //   7'h2F:
	        //     for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	        //       if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	        //         // Respective byte enables are asserted as per write strobes 
	        //         // Slave register 47
	        //         slv_reg47[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	        //       end  
	        //   7'h30:
	        //     for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	        //       if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	        //         // Respective byte enables are asserted as per write strobes 
	        //         // Slave register 48
	        //         slv_reg48[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	        //       end  
	        //   7'h31:
	        //     for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	        //       if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	        //         // Respective byte enables are asserted as per write strobes 
	        //         // Slave register 49
	        //         slv_reg49[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	        //       end  
	        //   7'h32:
	        //     for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	        //       if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	        //         // Respective byte enables are asserted as per write strobes 
	        //         // Slave register 50
	        //         slv_reg50[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	        //       end  
	        //   7'h33:
	        //     for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	        //       if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	        //         // Respective byte enables are asserted as per write strobes 
	        //         // Slave register 51
	        //         slv_reg51[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	        //       end  
	          7'h34:
	            for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	              if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	                // Respective byte enables are asserted as per write strobes 
	                // Slave register 52
	                slv_reg52[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	              end  
	          7'h35:
	            for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	              if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	                // Respective byte enables are asserted as per write strobes 
	                // Slave register 53
	                slv_reg53[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	              end  
	          7'h36:
	            for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	              if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	                // Respective byte enables are asserted as per write strobes 
	                // Slave register 54
	                slv_reg54[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	              end  
	          7'h37:
	            for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	              if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	                // Respective byte enables are asserted as per write strobes 
	                // Slave register 55
	                slv_reg55[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	              end  
	          7'h38:
	            for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	              if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	                // Respective byte enables are asserted as per write strobes 
	                // Slave register 56
	                slv_reg56[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	              end  
	          7'h39:
	            for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	              if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	                // Respective byte enables are asserted as per write strobes 
	                // Slave register 57
	                slv_reg57[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	              end  
	          7'h3A:
	            for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	              if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	                // Respective byte enables are asserted as per write strobes 
	                // Slave register 58
	                slv_reg58[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	              end  
	          7'h3B:
	            for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	              if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	                // Respective byte enables are asserted as per write strobes 
	                // Slave register 59
	                slv_reg59[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	              end  
	          7'h3C:
	            for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	              if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	                // Respective byte enables are asserted as per write strobes 
	                // Slave register 60
	                slv_reg60[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	              end  
	          7'h3D:
	            for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	              if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	                // Respective byte enables are asserted as per write strobes 
	                // Slave register 61
	                slv_reg61[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	              end  
	          7'h3E:
	            for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	              if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	                // Respective byte enables are asserted as per write strobes 
	                // Slave register 62
	                slv_reg62[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	              end  
	          7'h3F:
	            for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	              if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	                // Respective byte enables are asserted as per write strobes 
	                // Slave register 63
	                slv_reg63[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	              end  
	          default : begin
	                      slv_reg0 <= slv_reg0;
	                    //   slv_reg1 <= slv_reg1;
	                    //   slv_reg2 <= slv_reg2;
	                      slv_reg3 <= slv_reg3;
	                      slv_reg4 <= slv_reg4;
	                      slv_reg5 <= slv_reg5;
	                      slv_reg6 <= slv_reg6;
	                    //   slv_reg7 <= slv_reg7;
	                      slv_reg8 <= slv_reg8;
	                      slv_reg9 <= slv_reg9;
	                    //   slv_reg10 <= slv_reg10;
	                    //   slv_reg11 <= slv_reg11;
	                      slv_reg12 <= slv_reg12;
	                    //   slv_reg13 <= slv_reg13;
	                      slv_reg14 <= slv_reg14;
	                      slv_reg15 <= slv_reg15;
	                    //   slv_reg16 <= slv_reg16;
	                    //   slv_reg17 <= slv_reg17;
	                    //   slv_reg18 <= slv_reg18;
	                    //   slv_reg19 <= slv_reg19;
	                    //   slv_reg20 <= slv_reg20;
	                    //   slv_reg21 <= slv_reg21;
	                    //   slv_reg22 <= slv_reg22;
	                    //   slv_reg23 <= slv_reg23;
	                    //   slv_reg24 <= slv_reg24;
	                    //   slv_reg25 <= slv_reg25;
	                    //   slv_reg26 <= slv_reg26;
	                    //   slv_reg27 <= slv_reg27;
	                    //   slv_reg28 <= slv_reg28;
	                    //   slv_reg29 <= slv_reg29;
	                    //   slv_reg30 <= slv_reg30;
	                    //   slv_reg31 <= slv_reg31;
	                    //   slv_reg32 <= slv_reg32;
	                    //   slv_reg33 <= slv_reg33;
	                    //   slv_reg34 <= slv_reg34;
	                    //   slv_reg35 <= slv_reg35;
	                    //   slv_reg36 <= slv_reg36;
	                    //   slv_reg37 <= slv_reg37;
	                    //   slv_reg38 <= slv_reg38;
	                    //   slv_reg39 <= slv_reg39;
	                    //   slv_reg40 <= slv_reg40;
	                    //   slv_reg41 <= slv_reg41;
	                    //   slv_reg42 <= slv_reg42;
	                    //   slv_reg43 <= slv_reg43;
	                    //   slv_reg44 <= slv_reg44;
	                    //   slv_reg45 <= slv_reg45;
	                    //   slv_reg46 <= slv_reg46;
	                    //   slv_reg47 <= slv_reg47;
	                    //   slv_reg48 <= slv_reg48;
	                    //   slv_reg49 <= slv_reg49;
	                    //   slv_reg50 <= slv_reg50;
	                    //   slv_reg51 <= slv_reg51;
	                      slv_reg52 <= slv_reg52;
	                      slv_reg53 <= slv_reg53;
	                      slv_reg54 <= slv_reg54;
	                      slv_reg55 <= slv_reg55;
	                      slv_reg56 <= slv_reg56;
	                      slv_reg57 <= slv_reg57;
	                      slv_reg58 <= slv_reg58;
	                      slv_reg59 <= slv_reg59;
	                      slv_reg60 <= slv_reg60;
	                      slv_reg61 <= slv_reg61;
	                      slv_reg62 <= slv_reg62;
	                      slv_reg63 <= slv_reg63;
	                    end
	        endcase
	      end
	  end
	end   

	// Implement write response logic generation
	// The write response and response valid signals are asserted by the slave 
	// when axi_wready, S_AXI_WVALID, axi_wready and S_AXI_WVALID are asserted.  
	// This marks the acceptance of address and indicates the status of 
	// write transaction.

	always @( posedge S_AXI_ACLK )
	begin
	  if ( S_AXI_ARESETN == 1'b0 )
	    begin
	      axi_bvalid  <= 0;
	      axi_bresp   <= 2'b0;
	    end 
	  else
	    begin    
	      if (axi_awready && S_AXI_AWVALID && ~axi_bvalid && axi_wready && S_AXI_WVALID)
	        begin
	          // indicates a valid write response is available
	          axi_bvalid <= 1'b1;
	          axi_bresp  <= 2'b0; // 'OKAY' response 
	        end                   // work error responses in future
	      else
	        begin
	          if (S_AXI_BREADY && axi_bvalid) 
	            //check if bready is asserted while bvalid is high) 
	            //(there is a possibility that bready is always asserted high)   
	            begin
	              axi_bvalid <= 1'b0; 
	            end  
	        end
	    end
	end   

	// Implement axi_arready generation
	// axi_arready is asserted for one S_AXI_ACLK clock cycle when
	// S_AXI_ARVALID is asserted. axi_awready is 
	// de-asserted when reset (active low) is asserted. 
	// The read address is also latched when S_AXI_ARVALID is 
	// asserted. axi_araddr is reset to zero on reset assertion.

	always @( posedge S_AXI_ACLK )
	begin
	  if ( S_AXI_ARESETN == 1'b0 )
	    begin
	      axi_arready <= 1'b0;
	      axi_araddr  <= 32'b0;
	    end 
	  else
	    begin    
	      if (~axi_arready && S_AXI_ARVALID)
	        begin
	          // indicates that the slave has acceped the valid read address
	          axi_arready <= 1'b1;
	          // Read address latching
	          axi_araddr  <= S_AXI_ARADDR;
	        end
	      else
	        begin
	          axi_arready <= 1'b0;
	        end
	    end 
	end       

	// Implement axi_arvalid generation
	// axi_rvalid is asserted for one S_AXI_ACLK clock cycle when both 
	// S_AXI_ARVALID and axi_arready are asserted. The slave registers 
	// data are available on the axi_rdata bus at this instance. The 
	// assertion of axi_rvalid marks the validity of read data on the 
	// bus and axi_rresp indicates the status of read transaction.axi_rvalid 
	// is deasserted on reset (active low). axi_rresp and axi_rdata are 
	// cleared to zero on reset (active low).  
	always @( posedge S_AXI_ACLK )
	begin
	  if ( S_AXI_ARESETN == 1'b0 )
	    begin
	      axi_rvalid <= 0;
	      axi_rresp  <= 0;
	    end 
	  else
	    begin    
	      if (axi_arready && S_AXI_ARVALID && ~axi_rvalid)
	        begin
	          // Valid read data is available at the read data bus
	          axi_rvalid <= 1'b1;
	          axi_rresp  <= 2'b0; // 'OKAY' response
	        end   
	      else if (axi_rvalid && S_AXI_RREADY)
	        begin
	          // Read data is accepted by the master
	          axi_rvalid <= 1'b0;
	        end                
	    end
	end    

	// Implement memory mapped register select and read logic generation
	// Slave register read enable is asserted when valid address is available
	// and the slave is ready to accept the read address.
	assign slv_reg_rden = axi_arready & S_AXI_ARVALID & ~axi_rvalid;
	always @(*)
	begin
	      // Address decoding for reading registers
	      case ( axi_araddr[ADDR_LSB+OPT_MEM_ADDR_BITS:ADDR_LSB] )
	        7'h00   : reg_data_out <= slv_reg0;
	        7'h01   : reg_data_out <= slv_reg1;
	        7'h02   : reg_data_out <= slv_reg2;
	        7'h03   : reg_data_out <= slv_reg3;
	        7'h04   : reg_data_out <= slv_reg4;
	        7'h05   : reg_data_out <= slv_reg5;
	        7'h06   : reg_data_out <= slv_reg6;
	        7'h07   : reg_data_out <= slv_reg7;
	        7'h08   : reg_data_out <= slv_reg8;
	        7'h09   : reg_data_out <= slv_reg9;
	        7'h0A   : reg_data_out <= slv_reg10;
	        7'h0B   : reg_data_out <= slv_reg11;
	        7'h0C   : reg_data_out <= slv_reg12;
	        7'h0D   : reg_data_out <= slv_reg13;
	        7'h0E   : reg_data_out <= slv_reg14;
	        7'h0F   : reg_data_out <= slv_reg15;
	        7'h10   : reg_data_out <= slv_reg16;
	        7'h11   : reg_data_out <= slv_reg17;
	        7'h12   : reg_data_out <= slv_reg18;
	        7'h13   : reg_data_out <= slv_reg19;
	        7'h14   : reg_data_out <= slv_reg20;
	        7'h15   : reg_data_out <= slv_reg21;
	        7'h16   : reg_data_out <= slv_reg22;
	        7'h17   : reg_data_out <= slv_reg23;
	        7'h18   : reg_data_out <= slv_reg24;
	        7'h19   : reg_data_out <= slv_reg25;
	        7'h1A   : reg_data_out <= slv_reg26;
	        7'h1B   : reg_data_out <= slv_reg27;
	        7'h1C   : reg_data_out <= slv_reg28;
	        7'h1D   : reg_data_out <= slv_reg29;
	        7'h1E   : reg_data_out <= slv_reg30;
	        7'h1F   : reg_data_out <= slv_reg31;
	        7'h20   : reg_data_out <= slv_reg32;
	        7'h21   : reg_data_out <= slv_reg33;
	        7'h22   : reg_data_out <= slv_reg34;
	        7'h23   : reg_data_out <= slv_reg35;
	        7'h24   : reg_data_out <= slv_reg36;
	        7'h25   : reg_data_out <= slv_reg37;
	        7'h26   : reg_data_out <= slv_reg38;
	        7'h27   : reg_data_out <= slv_reg39;
	        7'h28   : reg_data_out <= slv_reg40;
	        7'h29   : reg_data_out <= slv_reg41;
	        7'h2A   : reg_data_out <= slv_reg42;
	        7'h2B   : reg_data_out <= slv_reg43;
	        7'h2C   : reg_data_out <= slv_reg44;
	        7'h2D   : reg_data_out <= slv_reg45;
	        7'h2E   : reg_data_out <= slv_reg46;
	        7'h2F   : reg_data_out <= slv_reg47;
	        7'h30   : reg_data_out <= slv_reg48;
	        7'h31   : reg_data_out <= slv_reg49;
	        7'h32   : reg_data_out <= slv_reg50;
	        7'h33   : reg_data_out <= slv_reg51;
	        7'h34   : reg_data_out <= slv_reg52;
	        7'h35   : reg_data_out <= slv_reg53;
	        7'h36   : reg_data_out <= slv_reg54;
	        7'h37   : reg_data_out <= slv_reg55;
	        7'h38   : reg_data_out <= slv_reg56;
	        7'h39   : reg_data_out <= slv_reg57;
	        7'h3A   : reg_data_out <= slv_reg58;
	        7'h3B   : reg_data_out <= slv_reg59;
	        7'h3C   : reg_data_out <= slv_reg60;
	        7'h3D   : reg_data_out <= slv_reg61;
	        7'h3E   : reg_data_out <= slv_reg62;
	        7'h3F   : reg_data_out <= slv_reg63;
	        default : reg_data_out <= 0;
	      endcase
	end

	// Output register or memory read data
	always @( posedge S_AXI_ACLK )
	begin
	  if ( S_AXI_ARESETN == 1'b0 )
	    begin
	      axi_rdata  <= 0;
	    end 
	  else
	    begin    
	      // When there is a valid read address (S_AXI_ARVALID) with 
	      // acceptance of read address by the slave (axi_arready), 
	      // output the read dada 
	      if (slv_reg_rden)
	        begin
	          axi_rdata <= reg_data_out;     // register read data
	        end   
	    end
	end    

	// Add user logic here

	// Write
	always @(posedge S_AXI_ACLK)
    begin
		o_WF_total_count		<= slv_reg0;
		o_WF_BRAM_WE			<= slv_reg3 [0];
		o_WF_start_count		<= slv_reg3 [1];
		o_WF_reset_count		<= slv_reg3 [2];
		o_WF_mode_sel			<= slv_reg3 [8];
		o_WF_addr				<= slv_reg4 [9:0];
		o_WF_data				<= slv_reg5;
		o_WF_dsp				<= slv_reg6 [15:0];
		o_c_factor				<= slv_reg8;
		o_v_factor				<= slv_reg9;
		o_Ready					<= slv_reg12 [0];
		o_Hart_beat				<= slv_reg12 [1];
		o_Write_Index			<= slv_reg60 [15:0];
		o_Write_DATA			<= slv_reg61;

		o_test_dpbram_addr		<= slv_reg62;
		o_test_dpbram_en		<= slv_reg63[0];
		o_test_dpbram_w_en		<= slv_reg63[1];
		o_test_dpbram_DSP_intr	<= slv_reg63[2];
		o_test_dpbram_wdata		<= slv_reg52;
		
    end

	// Read
	always @(posedge S_AXI_ACLK)
    begin
		slv_reg1 [0] 		<= i_WF_INT_0;
		slv_reg1 [1]		<= i_WF_INT_500;
		slv_reg2 			<= i_WF_current_count;
		slv_reg10			<= i_Float_ADC_C;
		slv_reg11			<= i_Float_ADC_V;
		slv_reg13 [0]		<= i_valid;
		slv_reg13 [1]		<= i_DSP_fail;
		slv_reg13 [2]		<= i_DSP_nENPWM;
		slv_reg16 			<= i_DSP_Duty;
		slv_reg17 [15:0] 	<= i_DSP_FaultNum;
		slv_reg18 			<= i_DSP_System_Status;
		slv_reg19 [15:0] 	<= i_DSP_EIS;
		slv_reg20 			<= i_DSP_RLoad;
		slv_reg21 [15:0] 	<= i_DSP_MPS_TYPE;
		slv_reg22 			<= i_DSP_SetCurrRD;
		slv_reg23 			<= i_DSP_DEGCurrentRD;
		slv_reg24 			<= i_DSP_DEGPeriod;
		slv_reg25 			<= i_DSP_OverCurrent;
		slv_reg26 			<= i_DSP_LowVoltage;
		slv_reg27 			<= i_DSP_OverVoltage;
		slv_reg28 			<= i_DSP_OverTemp;
		slv_reg29 			<= i_DSP_CurrentHighLimit;
		slv_reg30 			<= i_DSP_Vpgain;
		slv_reg31 			<= i_DSP_ViGain;
		slv_reg32 			<= i_DSP_CurrentPgain;
		slv_reg33 			<= i_DSP_CurrentIgain;
		slv_reg34 			<= i_DSP_Max_Duty;
		slv_reg35 [15:0] 	<= i_DSP_DSP_Code;
		slv_reg36 [15:0] 	<= i_DSP_SlewRate;
		slv_reg37 [15:0] 	<= i_DSP_osc_state;
		slv_reg38 [15:0] 	<= i_DSP_remote_state;
		slv_reg39 			<= i_DSP_regulation_time;
		slv_reg40 			<= i_DSP_Current_Factor;
		slv_reg41 			<= i_DSP_Voltage_Factor;
		slv_reg42 			<= i_DSP_Input_Voltage_Factor;
		slv_reg43 			<= i_DSP_Current_Offset_Set;
		slv_reg44 [15:0] 	<= i_DSP_Deadband_Set;
		slv_reg45 [15:0] 	<= i_DSP_Dual_Offset_Deadband_Set;
		slv_reg46 			<= i_DSP_PI_Max_V;
		slv_reg47 			<= i_DSP_PI_Min_V;
		slv_reg48 			<= i_DSP_Eruption_V;
		slv_reg49 			<= i_DSP_Eruption_C;
		slv_reg50 			<= i_F_DSP_ADC_C;
		slv_reg51 			<= i_F_DSP_ADC_V;

		slv_reg7			<= i_test_dpbram_rdata;
	end

	// User logic ends

endmodule